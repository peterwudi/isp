
module processing(
	input					clk,
	input		[31:0]	iData,



	output	[31:0]	oData
);



















endmodule
