// megafunction wizard: %Shift register (RAM-based)%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSHIFT_TAPS 

// ============================================================
// File Name: filter_shift_reg.v
// Megafunction Name(s):
// 			ALTSHIFT_TAPS
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module filter_shift_reg (
	clken,
	clock,
	shiftin,
	shiftout,
	taps0x,
	taps1x,
	taps2x);

	input	  clken;
	input	  clock;
	input	[23:0]  shiftin;
	output	[23:0]  shiftout;
	output	[23:0]  taps0x;
	output	[23:0]  taps1x;
	output	[23:0]  taps2x;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_off
`endif
	tri1	  clken;
`ifndef ALTERA_RESERVED_QIS
// synopsys translate_on
`endif

	wire [23:0] sub_wire0;
	wire [71:0] sub_wire1;
	wire [23:0] shiftout = sub_wire0[23:0];
	wire [47:24] sub_wire5 = sub_wire1[47:24];
	wire [71:48] sub_wire4 = sub_wire1[71:48];
	wire [71:48] sub_wire3 = sub_wire4[71:48];
	wire [23:0] sub_wire2 = sub_wire1[23:0];
	wire [23:0] taps0x = sub_wire2[23:0];
	wire [23:0] taps2x = sub_wire3[71:48];
	wire [23:0] taps1x = sub_wire5[47:24];

	altshift_taps	ALTSHIFT_TAPS_component (
				.clock (clock),
				.clken (clken),
				.shiftin (shiftin),
				.shiftout (sub_wire0),
				.taps (sub_wire1)
				// synopsys translate_off
				,
				.aclr ()
				// synopsys translate_on
				);
	defparam
		ALTSHIFT_TAPS_component.intended_device_family = "Stratix III",
		ALTSHIFT_TAPS_component.lpm_hint = "RAM_BLOCK_TYPE=AUTO",
		ALTSHIFT_TAPS_component.lpm_type = "altshift_taps",
		ALTSHIFT_TAPS_component.number_of_taps = 3,
		ALTSHIFT_TAPS_component.tap_distance = 322,
		ALTSHIFT_TAPS_component.width = 24;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: ACLR NUMERIC "0"
// Retrieval info: PRIVATE: CLKEN NUMERIC "1"
// Retrieval info: PRIVATE: GROUP_TAPS NUMERIC "1"
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: PRIVATE: NUMBER_OF_TAPS NUMERIC "3"
// Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "3"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: TAP_DISTANCE NUMERIC "322"
// Retrieval info: PRIVATE: WIDTH NUMERIC "24"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
// Retrieval info: CONSTANT: LPM_HINT STRING "RAM_BLOCK_TYPE=AUTO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "altshift_taps"
// Retrieval info: CONSTANT: NUMBER_OF_TAPS NUMERIC "3"
// Retrieval info: CONSTANT: TAP_DISTANCE NUMERIC "322"
// Retrieval info: CONSTANT: WIDTH NUMERIC "24"
// Retrieval info: USED_PORT: clken 0 0 0 0 INPUT VCC "clken"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: shiftin 0 0 24 0 INPUT NODEFVAL "shiftin[23..0]"
// Retrieval info: USED_PORT: shiftout 0 0 24 0 OUTPUT NODEFVAL "shiftout[23..0]"
// Retrieval info: USED_PORT: taps0x 0 0 24 0 OUTPUT NODEFVAL "taps0x[23..0]"
// Retrieval info: USED_PORT: taps1x 0 0 24 0 OUTPUT NODEFVAL "taps1x[23..0]"
// Retrieval info: USED_PORT: taps2x 0 0 24 0 OUTPUT NODEFVAL "taps2x[23..0]"
// Retrieval info: CONNECT: @clken 0 0 0 0 clken 0 0 0 0
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @shiftin 0 0 24 0 shiftin 0 0 24 0
// Retrieval info: CONNECT: shiftout 0 0 24 0 @shiftout 0 0 24 0
// Retrieval info: CONNECT: taps0x 0 0 24 0 @taps 0 0 24 0
// Retrieval info: CONNECT: taps1x 0 0 24 0 @taps 0 0 24 24
// Retrieval info: CONNECT: taps2x 0 0 24 0 @taps 0 0 24 48
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL filter_shift_reg_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
