module conveng
(
	input					clk,
	input					reset,

	input		[23:0]	iData,
	input					iValid,
	
	output				oReq,
	output	[23:0]	oData,
	output				oValid,
	output				oDone
);

parameter	width			= 1920;
parameter	height		= 1080;














endmodule
