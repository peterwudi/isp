



module isp (
	input					clk;
	

	output				out;
);









