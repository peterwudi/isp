// ddr2_sys.v

// Generated using ACDS version 13.0sp1 232 at 2013.10.25.16:21:32

`timescale 1 ps / 1 ps
module ddr2_sys (
		input  wire        clk_clk,          //    clk.clk
		input  wire        reset_reset_n,    //  reset.reset_n
		output wire [13:0] memory_mem_a,     // memory.mem_a
		output wire [1:0]  memory_mem_ba,    //       .mem_ba
		output wire [1:0]  memory_mem_ck,    //       .mem_ck
		output wire [1:0]  memory_mem_ck_n,  //       .mem_ck_n
		output wire [1:0]  memory_mem_cke,   //       .mem_cke
		output wire [1:0]  memory_mem_cs_n,  //       .mem_cs_n
		output wire [7:0]  memory_mem_dm,    //       .mem_dm
		output wire [0:0]  memory_mem_ras_n, //       .mem_ras_n
		output wire [0:0]  memory_mem_cas_n, //       .mem_cas_n
		output wire [0:0]  memory_mem_we_n,  //       .mem_we_n
		inout  wire [63:0] memory_mem_dq,    //       .mem_dq
		inout  wire [7:0]  memory_mem_dqs,   //       .mem_dqs
		inout  wire [7:0]  memory_mem_dqs_n, //       .mem_dqs_n
		output wire [1:0]  memory_mem_odt,   //       .mem_odt
		input  wire        oct_rdn,          //    oct.rdn
		input  wire        oct_rup           //       .rup
	);

	wire          ddr2_afi_clk_clk;                                                              // ddr2:afi_clk -> [crosser:out_clk, crosser_001:in_clk, ddr2_avl_translator:clk, ddr2_avl_translator_avalon_universal_slave_0_agent:clk, ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, rsp_xbar_demux:clk, rst_controller_002:clk, width_adapter:clk, width_adapter_001:clk]
	wire          master_0_master_waitrequest;                                                   // master_0_master_translator:av_waitrequest -> master_0:master_waitrequest
	wire   [31:0] master_0_master_writedata;                                                     // master_0:master_writedata -> master_0_master_translator:av_writedata
	wire   [31:0] master_0_master_address;                                                       // master_0:master_address -> master_0_master_translator:av_address
	wire          master_0_master_write;                                                         // master_0:master_write -> master_0_master_translator:av_write
	wire          master_0_master_read;                                                          // master_0:master_read -> master_0_master_translator:av_read
	wire   [31:0] master_0_master_readdata;                                                      // master_0_master_translator:av_readdata -> master_0:master_readdata
	wire    [3:0] master_0_master_byteenable;                                                    // master_0:master_byteenable -> master_0_master_translator:av_byteenable
	wire          master_0_master_readdatavalid;                                                 // master_0_master_translator:av_readdatavalid -> master_0:master_readdatavalid
	wire          ddr2_avl_translator_avalon_anti_slave_0_waitrequest;                           // ddr2:avl_ready -> ddr2_avl_translator:av_waitrequest
	wire    [2:0] ddr2_avl_translator_avalon_anti_slave_0_burstcount;                            // ddr2_avl_translator:av_burstcount -> ddr2:avl_size
	wire  [255:0] ddr2_avl_translator_avalon_anti_slave_0_writedata;                             // ddr2_avl_translator:av_writedata -> ddr2:avl_wdata
	wire   [24:0] ddr2_avl_translator_avalon_anti_slave_0_address;                               // ddr2_avl_translator:av_address -> ddr2:avl_addr
	wire          ddr2_avl_translator_avalon_anti_slave_0_write;                                 // ddr2_avl_translator:av_write -> ddr2:avl_write_req
	wire          ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer;                    // ddr2_avl_translator:av_beginbursttransfer -> ddr2:avl_burstbegin
	wire          ddr2_avl_translator_avalon_anti_slave_0_read;                                  // ddr2_avl_translator:av_read -> ddr2:avl_read_req
	wire  [255:0] ddr2_avl_translator_avalon_anti_slave_0_readdata;                              // ddr2:avl_rdata -> ddr2_avl_translator:av_readdata
	wire          ddr2_avl_translator_avalon_anti_slave_0_readdatavalid;                         // ddr2:avl_rdata_valid -> ddr2_avl_translator:av_readdatavalid
	wire   [31:0] ddr2_avl_translator_avalon_anti_slave_0_byteenable;                            // ddr2_avl_translator:av_byteenable -> ddr2:avl_be
	wire          master_0_master_translator_avalon_universal_master_0_waitrequest;              // master_0_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_0_master_translator:uav_waitrequest
	wire    [2:0] master_0_master_translator_avalon_universal_master_0_burstcount;               // master_0_master_translator:uav_burstcount -> master_0_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_writedata;                // master_0_master_translator:uav_writedata -> master_0_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_address;                  // master_0_master_translator:uav_address -> master_0_master_translator_avalon_universal_master_0_agent:av_address
	wire          master_0_master_translator_avalon_universal_master_0_lock;                     // master_0_master_translator:uav_lock -> master_0_master_translator_avalon_universal_master_0_agent:av_lock
	wire          master_0_master_translator_avalon_universal_master_0_write;                    // master_0_master_translator:uav_write -> master_0_master_translator_avalon_universal_master_0_agent:av_write
	wire          master_0_master_translator_avalon_universal_master_0_read;                     // master_0_master_translator:uav_read -> master_0_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] master_0_master_translator_avalon_universal_master_0_readdata;                 // master_0_master_translator_avalon_universal_master_0_agent:av_readdata -> master_0_master_translator:uav_readdata
	wire          master_0_master_translator_avalon_universal_master_0_debugaccess;              // master_0_master_translator:uav_debugaccess -> master_0_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] master_0_master_translator_avalon_universal_master_0_byteenable;               // master_0_master_translator:uav_byteenable -> master_0_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          master_0_master_translator_avalon_universal_master_0_readdatavalid;            // master_0_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_0_master_translator:uav_readdatavalid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // ddr2_avl_translator:uav_waitrequest -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [7:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;              // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_avl_translator:uav_burstcount
	wire  [255:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata;               // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_avl_translator:uav_writedata
	wire   [31:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address;                 // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_avl_translator:uav_address
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write;                   // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_avl_translator:uav_write
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock;                    // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_avl_translator:uav_lock
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read;                    // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_avl_translator:uav_read
	wire  [255:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                // ddr2_avl_translator:uav_readdata -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // ddr2_avl_translator:uav_readdatavalid -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_avl_translator:uav_debugaccess
	wire   [31:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;              // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_avl_translator:uav_byteenable
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;            // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [356:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data;             // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;            // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [356:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [257:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [257:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket;     // master_0_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_valid;           // master_0_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket;   // master_0_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [103:0] master_0_master_translator_avalon_universal_master_0_agent_cp_data;            // master_0_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          master_0_master_translator_avalon_universal_master_0_agent_cp_ready;           // addr_router:sink_ready -> master_0_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid;                   // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [355:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data;                    // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> ddr2:soft_reset_n
	wire          ddr2_afi_reset_reset;                                                          // ddr2:afi_reset_n -> [rst_controller:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                            // rst_controller_001:reset_out -> [addr_router:reset, cmd_xbar_demux:reset, crosser:in_reset, crosser_001:out_reset, master_0_master_translator:reset, master_0_master_translator_avalon_universal_master_0_agent:reset]
	wire          rst_controller_002_reset_out_reset;                                            // rst_controller_002:reset_out -> [crosser:out_reset, crosser_001:in_reset, ddr2_avl_translator:reset, ddr2_avl_translator_avalon_universal_slave_0_agent:reset, ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, rsp_xbar_demux:reset, width_adapter:reset, width_adapter_001:reset]
	wire          addr_router_src_endofpacket;                                                   // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                         // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                 // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [103:0] addr_router_src_data;                                                          // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [0:0] addr_router_src_channel;                                                       // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                         // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          crosser_001_out_ready;                                                         // master_0_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_001:out_ready
	wire          crosser_out_ready;                                                             // width_adapter:in_ready -> crosser:out_ready
	wire          width_adapter_src_endofpacket;                                                 // width_adapter:out_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_src_valid;                                                       // width_adapter:out_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_src_startofpacket;                                               // width_adapter:out_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [355:0] width_adapter_src_data;                                                        // width_adapter:out_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_src_ready;                                                       // ddr2_avl_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter:out_ready
	wire    [0:0] width_adapter_src_channel;                                                     // width_adapter:out_channel -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_src_endofpacket;                                                     // id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_src_valid;                                                           // id_router:src_valid -> width_adapter_001:in_valid
	wire          id_router_src_startofpacket;                                                   // id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [355:0] id_router_src_data;                                                            // id_router:src_data -> width_adapter_001:in_data
	wire    [0:0] id_router_src_channel;                                                         // id_router:src_channel -> width_adapter_001:in_channel
	wire          id_router_src_ready;                                                           // width_adapter_001:in_ready -> id_router:src_ready
	wire          width_adapter_001_src_endofpacket;                                             // width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                   // width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_001_src_startofpacket;                                           // width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [103:0] width_adapter_001_src_data;                                                    // width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	wire          width_adapter_001_src_ready;                                                   // rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	wire    [0:0] width_adapter_001_src_channel;                                                 // width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	wire          crosser_out_endofpacket;                                                       // crosser:out_endofpacket -> width_adapter:in_endofpacket
	wire          crosser_out_valid;                                                             // crosser:out_valid -> width_adapter:in_valid
	wire          crosser_out_startofpacket;                                                     // crosser:out_startofpacket -> width_adapter:in_startofpacket
	wire  [103:0] crosser_out_data;                                                              // crosser:out_data -> width_adapter:in_data
	wire          crosser_out_channel;                                                           // crosser:out_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src0_endofpacket;                                               // cmd_xbar_demux:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                     // cmd_xbar_demux:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                             // cmd_xbar_demux:src0_startofpacket -> crosser:in_startofpacket
	wire  [103:0] cmd_xbar_demux_src0_data;                                                      // cmd_xbar_demux:src0_data -> crosser:in_data
	wire    [0:0] cmd_xbar_demux_src0_channel;                                                   // cmd_xbar_demux:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                     // crosser:in_ready -> cmd_xbar_demux:src0_ready
	wire          crosser_001_out_endofpacket;                                                   // crosser_001:out_endofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_001_out_valid;                                                         // crosser_001:out_valid -> master_0_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_001_out_startofpacket;                                                 // crosser_001:out_startofpacket -> master_0_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [103:0] crosser_001_out_data;                                                          // crosser_001:out_data -> master_0_master_translator_avalon_universal_master_0_agent:rp_data
	wire          crosser_001_out_channel;                                                       // crosser_001:out_channel -> master_0_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                               // rsp_xbar_demux:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                     // rsp_xbar_demux:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                             // rsp_xbar_demux:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [103:0] rsp_xbar_demux_src0_data;                                                      // rsp_xbar_demux:src0_data -> crosser_001:in_data
	wire    [0:0] rsp_xbar_demux_src0_channel;                                                   // rsp_xbar_demux:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                     // crosser_001:in_ready -> rsp_xbar_demux:src0_ready

	ddr2_sys_ddr2 ddr2 (
		.pll_ref_clk        (clk_clk),                                                    //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                              //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_reset_out_reset),                            //       soft_reset.reset_n
		.afi_clk            (ddr2_afi_clk_clk),                                           //          afi_clk.clk
		.afi_half_clk       (),                                                           //     afi_half_clk.clk
		.afi_reset_n        (ddr2_afi_reset_reset),                                       //        afi_reset.reset_n
		.afi_reset_export_n (),                                                           // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                               //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                              //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                              //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                            //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                             //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                            //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                              //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                           //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                           //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                            //                 .mem_we_n
		.mem_dq             (memory_mem_dq),                                              //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                             //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                           //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                             //                 .mem_odt
		.avl_ready          (ddr2_avl_translator_avalon_anti_slave_0_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (ddr2_avl_translator_avalon_anti_slave_0_address),            //                 .address
		.avl_rdata_valid    (ddr2_avl_translator_avalon_anti_slave_0_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (ddr2_avl_translator_avalon_anti_slave_0_readdata),           //                 .readdata
		.avl_wdata          (ddr2_avl_translator_avalon_anti_slave_0_writedata),          //                 .writedata
		.avl_be             (ddr2_avl_translator_avalon_anti_slave_0_byteenable),         //                 .byteenable
		.avl_read_req       (ddr2_avl_translator_avalon_anti_slave_0_read),               //                 .read
		.avl_write_req      (ddr2_avl_translator_avalon_anti_slave_0_write),              //                 .write
		.avl_size           (ddr2_avl_translator_avalon_anti_slave_0_burstcount),         //                 .burstcount
		.local_init_done    (),                                                           //           status.local_init_done
		.local_cal_success  (),                                                           //                 .local_cal_success
		.local_cal_fail     (),                                                           //                 .local_cal_fail
		.oct_rdn            (oct_rdn),                                                    //              oct.rdn
		.oct_rup            (oct_rup)                                                     //                 .rup
	);

	ddr2_sys_master_0 #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_0 (
		.clk_clk              (clk_clk),                       //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                //    clk_reset.reset
		.master_address       (master_0_master_address),       //       master.address
		.master_readdata      (master_0_master_readdata),      //             .readdata
		.master_read          (master_0_master_read),          //             .read
		.master_write         (master_0_master_write),         //             .write
		.master_writedata     (master_0_master_writedata),     //             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                               // master_reset.reset
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_0_master_translator (
		.clk                      (clk_clk),                                                            //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                 //                     reset.reset
		.uav_address              (master_0_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (master_0_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (master_0_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (master_0_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (master_0_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (master_0_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (master_0_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (master_0_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (master_0_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (master_0_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (master_0_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (master_0_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (master_0_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (master_0_master_byteenable),                                         //                          .byteenable
		.av_read                  (master_0_master_read),                                               //                          .read
		.av_readdata              (master_0_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (master_0_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (master_0_master_write),                                              //                          .write
		.av_writedata             (master_0_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.av_debugaccess           (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (256),
		.UAV_DATA_W                     (256),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (32),
		.UAV_BYTEENABLE_W               (32),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (8),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (32),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_avl_translator (
		.clk                      (ddr2_afi_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (ddr2_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~ddr2_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (97),
		.PKT_PROTECTION_L          (95),
		.PKT_BEGIN_BURST           (90),
		.PKT_BURSTWRAP_H           (82),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (85),
		.PKT_BURST_SIZE_L          (83),
		.PKT_BURST_TYPE_H          (87),
		.PKT_BURST_TYPE_L          (86),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (92),
		.PKT_SRC_ID_L              (92),
		.PKT_DEST_ID_H             (93),
		.PKT_DEST_ID_L             (93),
		.PKT_THREAD_ID_H           (94),
		.PKT_THREAD_ID_L           (94),
		.PKT_CACHE_H               (101),
		.PKT_CACHE_L               (98),
		.PKT_DATA_SIDEBAND_H       (89),
		.PKT_DATA_SIDEBAND_L       (89),
		.PKT_QOS_H                 (91),
		.PKT_QOS_L                 (91),
		.PKT_ADDR_SIDEBAND_H       (88),
		.PKT_ADDR_SIDEBAND_L       (88),
		.PKT_RESPONSE_STATUS_H     (103),
		.PKT_RESPONSE_STATUS_L     (102),
		.ST_DATA_W                 (104),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) master_0_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                     //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.av_address              (master_0_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (master_0_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (master_0_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (master_0_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (master_0_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (master_0_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (master_0_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (master_0_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (master_0_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (master_0_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (master_0_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (crosser_001_out_valid),                                                       //        rp.valid
		.rp_data                 (crosser_001_out_data),                                                        //          .data
		.rp_channel              (crosser_001_out_channel),                                                     //          .channel
		.rp_startofpacket        (crosser_001_out_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (crosser_001_out_endofpacket),                                                 //          .endofpacket
		.rp_ready                (crosser_001_out_ready),                                                       //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (342),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_ADDR_H                (319),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (320),
		.PKT_TRANS_POSTED          (321),
		.PKT_TRANS_WRITE           (322),
		.PKT_TRANS_READ            (323),
		.PKT_TRANS_LOCK            (324),
		.PKT_SRC_ID_H              (344),
		.PKT_SRC_ID_L              (344),
		.PKT_DEST_ID_H             (345),
		.PKT_DEST_ID_L             (345),
		.PKT_BURSTWRAP_H           (334),
		.PKT_BURSTWRAP_L           (334),
		.PKT_BYTE_CNT_H            (333),
		.PKT_BYTE_CNT_L            (326),
		.PKT_PROTECTION_H          (349),
		.PKT_PROTECTION_L          (347),
		.PKT_RESPONSE_STATUS_H     (355),
		.PKT_RESPONSE_STATUS_L     (354),
		.PKT_BURST_SIZE_H          (337),
		.PKT_BURST_SIZE_L          (335),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (356),
		.AVS_BURSTCOUNT_W          (8),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_src_ready),                                                       //              cp.ready
		.cp_valid                (width_adapter_src_valid),                                                       //                .valid
		.cp_data                 (width_adapter_src_data),                                                        //                .data
		.cp_startofpacket        (width_adapter_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (width_adapter_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (width_adapter_src_channel),                                                     //                .channel
		.rf_sink_ready           (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (357),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (258),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (ddr2_afi_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                      // clk_reset.reset
		.in_data           (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	ddr2_sys_addr_router addr_router (
		.sink_ready         (master_0_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (master_0_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (master_0_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (master_0_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (master_0_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_src_valid),                                                       //          .valid
		.src_data           (addr_router_src_data),                                                        //          .data
		.src_channel        (addr_router_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                  //          .endofpacket
	);

	ddr2_sys_id_router id_router (
		.sink_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_afi_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                 //       src.ready
		.src_valid          (id_router_src_valid),                                                 //          .valid
		.src_data           (id_router_src_data),                                                  //          .data
		.src_channel        (id_router_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                            //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.reset_in1  (~ddr2_afi_reset_reset),          // reset_in1.reset
		.clk        (),                               //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~ddr2_afi_reset_reset),              // reset_in0.reset
		.clk        (ddr2_afi_clk_clk),                   //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	ddr2_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                            //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	ddr2_sys_cmd_xbar_demux rsp_xbar_demux (
		.clk                (ddr2_afi_clk_clk),                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),       //          .channel
		.sink_data          (width_adapter_001_src_data),          //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),           //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),           //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),            //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),         //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),   //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)      //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (82),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (85),
		.IN_PKT_BURST_SIZE_L           (83),
		.IN_PKT_RESPONSE_STATUS_H      (103),
		.IN_PKT_RESPONSE_STATUS_L      (102),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (87),
		.IN_PKT_BURST_TYPE_L           (86),
		.IN_ST_DATA_W                  (104),
		.OUT_PKT_ADDR_H                (319),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (333),
		.OUT_PKT_BYTE_CNT_L            (326),
		.OUT_PKT_TRANS_COMPRESSED_READ (320),
		.OUT_PKT_BURST_SIZE_H          (337),
		.OUT_PKT_BURST_SIZE_L          (335),
		.OUT_PKT_RESPONSE_STATUS_H     (355),
		.OUT_PKT_RESPONSE_STATUS_L     (354),
		.OUT_PKT_TRANS_EXCLUSIVE       (325),
		.OUT_PKT_BURST_TYPE_H          (339),
		.OUT_PKT_BURST_TYPE_L          (338),
		.OUT_ST_DATA_W                 (356),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (ddr2_afi_clk_clk),                   //       clk.clk
		.reset                (rst_controller_002_reset_out_reset), // clk_reset.reset
		.in_valid             (crosser_out_valid),                  //      sink.valid
		.in_channel           (crosser_out_channel),                //          .channel
		.in_startofpacket     (crosser_out_startofpacket),          //          .startofpacket
		.in_endofpacket       (crosser_out_endofpacket),            //          .endofpacket
		.in_ready             (crosser_out_ready),                  //          .ready
		.in_data              (crosser_out_data),                   //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (319),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (333),
		.IN_PKT_BYTE_CNT_L             (326),
		.IN_PKT_TRANS_COMPRESSED_READ  (320),
		.IN_PKT_BURSTWRAP_H            (334),
		.IN_PKT_BURSTWRAP_L            (334),
		.IN_PKT_BURST_SIZE_H           (337),
		.IN_PKT_BURST_SIZE_L           (335),
		.IN_PKT_RESPONSE_STATUS_H      (355),
		.IN_PKT_RESPONSE_STATUS_L      (354),
		.IN_PKT_TRANS_EXCLUSIVE        (325),
		.IN_PKT_BURST_TYPE_H           (339),
		.IN_PKT_BURST_TYPE_L           (338),
		.IN_ST_DATA_W                  (356),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (81),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (85),
		.OUT_PKT_BURST_SIZE_L          (83),
		.OUT_PKT_RESPONSE_STATUS_H     (103),
		.OUT_PKT_RESPONSE_STATUS_L     (102),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (87),
		.OUT_PKT_BURST_TYPE_L          (86),
		.OUT_ST_DATA_W                 (104),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (ddr2_afi_clk_clk),                    //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_src_valid),                 //      sink.valid
		.in_channel           (id_router_src_channel),               //          .channel
		.in_startofpacket     (id_router_src_startofpacket),         //          .startofpacket
		.in_endofpacket       (id_router_src_endofpacket),           //          .endofpacket
		.in_ready             (id_router_src_ready),                 //          .ready
		.in_data              (id_router_src_data),                  //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (104),
		.BITS_PER_SYMBOL     (104),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                            //        in_clk.clk
		.in_reset          (rst_controller_001_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (ddr2_afi_clk_clk),                   //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset), // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src0_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (104),
		.BITS_PER_SYMBOL     (104),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (1),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (ddr2_afi_clk_clk),                   //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (clk_clk),                            //       out_clk.clk
		.out_reset         (rst_controller_001_reset_out_reset), // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src0_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

endmodule
