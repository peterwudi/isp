// ddr2_sys.v

// Generated using ACDS version 13.0sp1 232 at 2013.10.26.15:45:45

`timescale 1 ps / 1 ps
module ddr2_sys (
		input  wire        clk_clk,                    //    clk.clk
		input  wire        reset_reset_n,              //  reset.reset_n
		output wire [13:0] memory_mem_a,               // memory.mem_a
		output wire [1:0]  memory_mem_ba,              //       .mem_ba
		output wire [1:0]  memory_mem_ck,              //       .mem_ck
		output wire [1:0]  memory_mem_ck_n,            //       .mem_ck_n
		output wire [1:0]  memory_mem_cke,             //       .mem_cke
		output wire [1:0]  memory_mem_cs_n,            //       .mem_cs_n
		output wire [7:0]  memory_mem_dm,              //       .mem_dm
		output wire [0:0]  memory_mem_ras_n,           //       .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,           //       .mem_cas_n
		output wire [0:0]  memory_mem_we_n,            //       .mem_we_n
		inout  wire [63:0] memory_mem_dq,              //       .mem_dq
		inout  wire [7:0]  memory_mem_dqs,             //       .mem_dqs
		inout  wire [7:0]  memory_mem_dqs_n,           //       .mem_dqs_n
		output wire [1:0]  memory_mem_odt,             //       .mem_odt
		input  wire        oct_rdn,                    //    oct.rdn
		input  wire        oct_rup,                    //       .rup
		input  wire [29:0] read_control_read_base,     //   read.control_read_base
		input  wire [29:0] read_control_read_length,   //       .control_read_length
		input  wire        read_control_go,            //       .control_go
		output wire        read_control_done,          //       .control_done
		output wire        read_control_early_done,    //       .control_early_done
		input  wire        read_user_read_buffer,      //       .user_read_buffer
		input  wire [31:0] read_user_buffer_data,      //       .user_buffer_data
		output wire        read_user_data_available,   //       .user_data_available
		input  wire [29:0] write_control_write_base,   //  write.control_write_base
		input  wire [29:0] write_control_write_length, //       .control_write_length
		input  wire        write_control_go,           //       .control_go
		output wire        write_control_done,         //       .control_done
		input  wire        write_user_write_buffer,    //       .user_write_buffer
		input  wire [31:0] write_user_buffer_data,     //       .user_buffer_data
		output wire        write_user_buffer_full      //       .user_buffer_full
	);

	wire          ddr2_afi_clk_clk;                                                               // ddr2:afi_clk -> [addr_router:clk, cmd_xbar_demux:clk, ddr2_avl_translator:clk, ddr2_avl_translator_avalon_universal_slave_0_agent:clk, ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, read:clk, read_avalon_master_translator:clk, read_avalon_master_translator_avalon_universal_master_0_agent:clk, rsp_xbar_demux:clk, rst_controller_001:clk, rst_controller_002:clk, width_adapter:clk, width_adapter_001:clk, write:clk]
	wire          read_avalon_master_waitrequest;                                                 // read_avalon_master_translator:av_waitrequest -> read:master_waitrequest
	wire   [29:0] read_avalon_master_address;                                                     // read:master_address -> read_avalon_master_translator:av_address
	wire          read_avalon_master_read;                                                        // read:master_read -> read_avalon_master_translator:av_read
	wire   [31:0] read_avalon_master_readdata;                                                    // read_avalon_master_translator:av_readdata -> read:master_readdata
	wire          read_avalon_master_readdatavalid;                                               // read_avalon_master_translator:av_readdatavalid -> read:master_readdatavalid
	wire    [3:0] read_avalon_master_byteenable;                                                  // read:master_byteenable -> read_avalon_master_translator:av_byteenable
	wire          ddr2_avl_translator_avalon_anti_slave_0_waitrequest;                            // ddr2:avl_ready -> ddr2_avl_translator:av_waitrequest
	wire    [2:0] ddr2_avl_translator_avalon_anti_slave_0_burstcount;                             // ddr2_avl_translator:av_burstcount -> ddr2:avl_size
	wire  [255:0] ddr2_avl_translator_avalon_anti_slave_0_writedata;                              // ddr2_avl_translator:av_writedata -> ddr2:avl_wdata
	wire   [24:0] ddr2_avl_translator_avalon_anti_slave_0_address;                                // ddr2_avl_translator:av_address -> ddr2:avl_addr
	wire          ddr2_avl_translator_avalon_anti_slave_0_write;                                  // ddr2_avl_translator:av_write -> ddr2:avl_write_req
	wire          ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer;                     // ddr2_avl_translator:av_beginbursttransfer -> ddr2:avl_burstbegin
	wire          ddr2_avl_translator_avalon_anti_slave_0_read;                                   // ddr2_avl_translator:av_read -> ddr2:avl_read_req
	wire  [255:0] ddr2_avl_translator_avalon_anti_slave_0_readdata;                               // ddr2:avl_rdata -> ddr2_avl_translator:av_readdata
	wire          ddr2_avl_translator_avalon_anti_slave_0_readdatavalid;                          // ddr2:avl_rdata_valid -> ddr2_avl_translator:av_readdatavalid
	wire   [31:0] ddr2_avl_translator_avalon_anti_slave_0_byteenable;                             // ddr2_avl_translator:av_byteenable -> ddr2:avl_be
	wire          read_avalon_master_translator_avalon_universal_master_0_waitrequest;            // read_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> read_avalon_master_translator:uav_waitrequest
	wire    [2:0] read_avalon_master_translator_avalon_universal_master_0_burstcount;             // read_avalon_master_translator:uav_burstcount -> read_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] read_avalon_master_translator_avalon_universal_master_0_writedata;              // read_avalon_master_translator:uav_writedata -> read_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [29:0] read_avalon_master_translator_avalon_universal_master_0_address;                // read_avalon_master_translator:uav_address -> read_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          read_avalon_master_translator_avalon_universal_master_0_lock;                   // read_avalon_master_translator:uav_lock -> read_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          read_avalon_master_translator_avalon_universal_master_0_write;                  // read_avalon_master_translator:uav_write -> read_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          read_avalon_master_translator_avalon_universal_master_0_read;                   // read_avalon_master_translator:uav_read -> read_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] read_avalon_master_translator_avalon_universal_master_0_readdata;               // read_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> read_avalon_master_translator:uav_readdata
	wire          read_avalon_master_translator_avalon_universal_master_0_debugaccess;            // read_avalon_master_translator:uav_debugaccess -> read_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] read_avalon_master_translator_avalon_universal_master_0_byteenable;             // read_avalon_master_translator:uav_byteenable -> read_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          read_avalon_master_translator_avalon_universal_master_0_readdatavalid;          // read_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> read_avalon_master_translator:uav_readdatavalid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // ddr2_avl_translator:uav_waitrequest -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [7:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount;               // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_avl_translator:uav_burstcount
	wire  [255:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata;                // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_avl_translator:uav_writedata
	wire   [29:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address;                  // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_avl_translator:uav_address
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write;                    // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_avl_translator:uav_write
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock;                     // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_avl_translator:uav_lock
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read;                     // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_avl_translator:uav_read
	wire  [255:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata;                 // ddr2_avl_translator:uav_readdata -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // ddr2_avl_translator:uav_readdatavalid -> ddr2_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_avl_translator:uav_debugaccess
	wire   [31:0] ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable;               // ddr2_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_avl_translator:uav_byteenable
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid;             // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [354:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data;              // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready;             // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [354:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // ddr2_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [257:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          read_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;   // read_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          read_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;         // read_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          read_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket; // read_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [101:0] read_avalon_master_translator_avalon_universal_master_0_agent_cp_data;          // read_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          read_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;         // addr_router:sink_ready -> read_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid;                    // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [353:0] ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data;                     // ddr2_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router:sink_ready -> ddr2_avl_translator_avalon_universal_slave_0_agent:rp_ready
	wire          rst_controller_reset_out_reset;                                                 // rst_controller:reset_out -> ddr2:soft_reset_n
	wire          ddr2_afi_reset_reset;                                                           // ddr2:afi_reset_n -> [rst_controller:reset_in1, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                                             // rst_controller_001:reset_out -> [addr_router:reset, cmd_xbar_demux:reset, read:reset, read_avalon_master_translator:reset, read_avalon_master_translator_avalon_universal_master_0_agent:reset, write:reset]
	wire          rst_controller_002_reset_out_reset;                                             // rst_controller_002:reset_out -> [ddr2_avl_translator:reset, ddr2_avl_translator_avalon_universal_slave_0_agent:reset, ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, rsp_xbar_demux:reset, width_adapter:reset, width_adapter_001:reset]
	wire          cmd_xbar_demux_src0_endofpacket;                                                // cmd_xbar_demux:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                      // cmd_xbar_demux:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                              // cmd_xbar_demux:src0_startofpacket -> width_adapter:in_startofpacket
	wire  [101:0] cmd_xbar_demux_src0_data;                                                       // cmd_xbar_demux:src0_data -> width_adapter:in_data
	wire    [0:0] cmd_xbar_demux_src0_channel;                                                    // cmd_xbar_demux:src0_channel -> width_adapter:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                // rsp_xbar_demux:src0_endofpacket -> read_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                      // rsp_xbar_demux:src0_valid -> read_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                              // rsp_xbar_demux:src0_startofpacket -> read_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [101:0] rsp_xbar_demux_src0_data;                                                       // rsp_xbar_demux:src0_data -> read_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_src0_channel;                                                    // rsp_xbar_demux:src0_channel -> read_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_src_endofpacket;                                                    // addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          addr_router_src_valid;                                                          // addr_router:src_valid -> cmd_xbar_demux:sink_valid
	wire          addr_router_src_startofpacket;                                                  // addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [101:0] addr_router_src_data;                                                           // addr_router:src_data -> cmd_xbar_demux:sink_data
	wire    [0:0] addr_router_src_channel;                                                        // addr_router:src_channel -> cmd_xbar_demux:sink_channel
	wire          addr_router_src_ready;                                                          // cmd_xbar_demux:sink_ready -> addr_router:src_ready
	wire          rsp_xbar_demux_src0_ready;                                                      // read_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux:src0_ready
	wire          cmd_xbar_demux_src0_ready;                                                      // width_adapter:in_ready -> cmd_xbar_demux:src0_ready
	wire          width_adapter_src_endofpacket;                                                  // width_adapter:out_endofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_src_valid;                                                        // width_adapter:out_valid -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_src_startofpacket;                                                // width_adapter:out_startofpacket -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [353:0] width_adapter_src_data;                                                         // width_adapter:out_data -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_src_ready;                                                        // ddr2_avl_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter:out_ready
	wire    [0:0] width_adapter_src_channel;                                                      // width_adapter:out_channel -> ddr2_avl_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_src_endofpacket;                                                      // id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_src_valid;                                                            // id_router:src_valid -> width_adapter_001:in_valid
	wire          id_router_src_startofpacket;                                                    // id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [353:0] id_router_src_data;                                                             // id_router:src_data -> width_adapter_001:in_data
	wire    [0:0] id_router_src_channel;                                                          // id_router:src_channel -> width_adapter_001:in_channel
	wire          id_router_src_ready;                                                            // width_adapter_001:in_ready -> id_router:src_ready
	wire          width_adapter_001_src_endofpacket;                                              // width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                    // width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_001_src_startofpacket;                                            // width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [101:0] width_adapter_001_src_data;                                                     // width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	wire          width_adapter_001_src_ready;                                                    // rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	wire    [0:0] width_adapter_001_src_channel;                                                  // width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel

	ddr2_sys_ddr2 ddr2 (
		.pll_ref_clk        (clk_clk),                                                    //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                              //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_reset_out_reset),                            //       soft_reset.reset_n
		.afi_clk            (ddr2_afi_clk_clk),                                           //          afi_clk.clk
		.afi_half_clk       (),                                                           //     afi_half_clk.clk
		.afi_reset_n        (ddr2_afi_reset_reset),                                       //        afi_reset.reset_n
		.afi_reset_export_n (),                                                           // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                               //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                              //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                              //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                            //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                             //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                            //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                              //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                           //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                           //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                            //                 .mem_we_n
		.mem_dq             (memory_mem_dq),                                              //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                             //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                           //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                             //                 .mem_odt
		.avl_ready          (ddr2_avl_translator_avalon_anti_slave_0_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (ddr2_avl_translator_avalon_anti_slave_0_address),            //                 .address
		.avl_rdata_valid    (ddr2_avl_translator_avalon_anti_slave_0_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (ddr2_avl_translator_avalon_anti_slave_0_readdata),           //                 .readdata
		.avl_wdata          (ddr2_avl_translator_avalon_anti_slave_0_writedata),          //                 .writedata
		.avl_be             (ddr2_avl_translator_avalon_anti_slave_0_byteenable),         //                 .byteenable
		.avl_read_req       (ddr2_avl_translator_avalon_anti_slave_0_read),               //                 .read
		.avl_write_req      (ddr2_avl_translator_avalon_anti_slave_0_write),              //                 .write
		.avl_size           (ddr2_avl_translator_avalon_anti_slave_0_burstcount),         //                 .burstcount
		.local_init_done    (),                                                           //           status.local_init_done
		.local_cal_success  (),                                                           //                 .local_cal_success
		.local_cal_fail     (),                                                           //                 .local_cal_fail
		.oct_rdn            (oct_rdn),                                                    //              oct.rdn
		.oct_rup            (oct_rup)                                                     //                 .rup
	);

	mem_read_buffer_avalon_interface #(
		.DATAWIDTH       (32),
		.BYTEENABLEWIDTH (4),
		.ADDRESSWIDTH    (30),
		.FIFODEPTH       (32),
		.FIFODEPTH_LOG2  (5),
		.FIFOUSEMEMORY   (1)
	) read (
		.reset                (rst_controller_001_reset_out_reset), //    reset_sink.reset
		.clk                  (ddr2_afi_clk_clk),                   //    clock_sink.clk
		.master_address       (read_avalon_master_address),         // avalon_master.address
		.master_read          (read_avalon_master_read),            //              .read
		.master_byteenable    (read_avalon_master_byteenable),      //              .byteenable
		.master_readdata      (read_avalon_master_readdata),        //              .readdata
		.master_readdatavalid (read_avalon_master_readdatavalid),   //              .readdatavalid
		.master_waitrequest   (read_avalon_master_waitrequest),     //              .waitrequest
		.control_read_base    (read_control_read_base),             //   conduit_end.export
		.control_read_length  (read_control_read_length),           //              .export
		.control_go           (read_control_go),                    //              .export
		.control_done         (read_control_done),                  //              .export
		.control_early_done   (read_control_early_done),            //              .export
		.user_read_buffer     (read_user_read_buffer),              //              .export
		.user_buffer_data     (read_user_buffer_data),              //              .export
		.user_data_available  (read_user_data_available)            //              .export
	);

	mem_write_buffer_avalon_interface #(
		.DATAWIDTH       (32),
		.BYTEENABLEWIDTH (4),
		.ADDRESSWIDTH    (30),
		.FIFODEPTH       (32),
		.FIFODEPTH_LOG2  (5),
		.FIFOUSEMEMORY   (1)
	) write (
		.clk                  (ddr2_afi_clk_clk),                   //    clock_sink.clk
		.reset                (rst_controller_001_reset_out_reset), //    reset_sink.reset
		.control_write_base   (write_control_write_base),           //   conduit_end.export
		.control_write_length (write_control_write_length),         //              .export
		.control_go           (write_control_go),                   //              .export
		.control_done         (write_control_done),                 //              .export
		.user_write_buffer    (write_user_write_buffer),            //              .export
		.user_buffer_data     (write_user_buffer_data),             //              .export
		.user_buffer_full     (write_user_buffer_full),             //              .export
		.master_address       (),                                   // avalon_master.address
		.master_write         (),                                   //              .write
		.master_byteenable    (),                                   //              .byteenable
		.master_writedata     (),                                   //              .writedata
		.master_waitrequest   ()                                    //              .waitrequest
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (30),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) read_avalon_master_translator (
		.clk                      (ddr2_afi_clk_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                    //                     reset.reset
		.uav_address              (read_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (read_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (read_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (read_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (read_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (read_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (read_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (read_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (read_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (read_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (read_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (read_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (read_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (read_avalon_master_byteenable),                                         //                          .byteenable
		.av_read                  (read_avalon_master_read),                                               //                          .read
		.av_readdata              (read_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (read_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_chipselect            (1'b0),                                                                  //               (terminated)
		.av_write                 (1'b0),                                                                  //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                  //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (256),
		.UAV_DATA_W                     (256),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (32),
		.UAV_BYTEENABLE_W               (32),
		.UAV_ADDRESS_W                  (30),
		.UAV_BURSTCOUNT_W               (8),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (32),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_avl_translator (
		.clk                      (ddr2_afi_clk_clk),                                                    //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                  //                    reset.reset
		.uav_address              (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_avl_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_avl_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_avl_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_avl_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_avl_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (ddr2_avl_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (ddr2_avl_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_avl_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_avl_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~ddr2_avl_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_chipselect            (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (72),
		.PKT_ADDR_H                (65),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (66),
		.PKT_TRANS_POSTED          (67),
		.PKT_TRANS_WRITE           (68),
		.PKT_TRANS_READ            (69),
		.PKT_TRANS_LOCK            (70),
		.PKT_TRANS_EXCLUSIVE       (71),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (92),
		.PKT_THREAD_ID_L           (92),
		.PKT_CACHE_H               (99),
		.PKT_CACHE_L               (96),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) read_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (ddr2_afi_clk_clk),                                                               //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.av_address              (read_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (read_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (read_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (read_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (read_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (read_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (read_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (read_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (read_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (read_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (read_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (read_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (read_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (read_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (read_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (read_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_src0_valid),                                                      //        rp.valid
		.rp_data                 (rsp_xbar_demux_src0_data),                                                       //          .data
		.rp_channel              (rsp_xbar_demux_src0_channel),                                                    //          .channel
		.rp_startofpacket        (rsp_xbar_demux_src0_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_src0_endofpacket),                                                //          .endofpacket
		.rp_ready                (rsp_xbar_demux_src0_ready),                                                      //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (255),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (340),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (287),
		.PKT_BYTEEN_L              (256),
		.PKT_ADDR_H                (317),
		.PKT_ADDR_L                (288),
		.PKT_TRANS_COMPRESSED_READ (318),
		.PKT_TRANS_POSTED          (319),
		.PKT_TRANS_WRITE           (320),
		.PKT_TRANS_READ            (321),
		.PKT_TRANS_LOCK            (322),
		.PKT_SRC_ID_H              (342),
		.PKT_SRC_ID_L              (342),
		.PKT_DEST_ID_H             (343),
		.PKT_DEST_ID_L             (343),
		.PKT_BURSTWRAP_H           (332),
		.PKT_BURSTWRAP_L           (332),
		.PKT_BYTE_CNT_H            (331),
		.PKT_BYTE_CNT_L            (324),
		.PKT_PROTECTION_H          (347),
		.PKT_PROTECTION_L          (345),
		.PKT_RESPONSE_STATUS_H     (353),
		.PKT_RESPONSE_STATUS_L     (352),
		.PKT_BURST_SIZE_H          (335),
		.PKT_BURST_SIZE_L          (333),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (354),
		.AVS_BURSTCOUNT_W          (8),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_avl_translator_avalon_universal_slave_0_agent (
		.clk                     (ddr2_afi_clk_clk),                                                              //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_avl_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_src_ready),                                                       //              cp.ready
		.cp_valid                (width_adapter_src_valid),                                                       //                .valid
		.cp_data                 (width_adapter_src_data),                                                        //                .data
		.cp_startofpacket        (width_adapter_src_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (width_adapter_src_endofpacket),                                                 //                .endofpacket
		.cp_channel              (width_adapter_src_channel),                                                     //                .channel
		.rf_sink_ready           (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (355),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (ddr2_afi_clk_clk),                                                              //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                            // clk_reset.reset
		.in_data           (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	ddr2_sys_addr_router addr_router (
		.sink_ready         (read_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (read_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (read_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (read_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (read_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (ddr2_afi_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_src_valid),                                                          //          .valid
		.src_data           (addr_router_src_data),                                                           //          .data
		.src_channel        (addr_router_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                     //          .endofpacket
	);

	ddr2_sys_id_router id_router (
		.sink_ready         (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (ddr2_afi_clk_clk),                                                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                 //       src.ready
		.src_valid          (id_router_src_valid),                                                 //          .valid
		.src_data           (id_router_src_data),                                                  //          .data
		.src_channel        (id_router_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                            //          .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (2),
		.OUTPUT_RESET_SYNC_EDGES ("none"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.reset_in1  (~ddr2_afi_reset_reset),          // reset_in1.reset
		.clk        (),                               //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (ddr2_afi_clk_clk),                   //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~ddr2_afi_reset_reset),              // reset_in0.reset
		.clk        (ddr2_afi_clk_clk),                   //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	ddr2_sys_cmd_xbar_demux cmd_xbar_demux (
		.clk                (ddr2_afi_clk_clk),                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sink_ready         (addr_router_src_ready),              //      sink.ready
		.sink_channel       (addr_router_src_channel),            //          .channel
		.sink_data          (addr_router_src_data),               //          .data
		.sink_startofpacket (addr_router_src_startofpacket),      //          .startofpacket
		.sink_endofpacket   (addr_router_src_endofpacket),        //          .endofpacket
		.sink_valid         (addr_router_src_valid),              //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	ddr2_sys_cmd_xbar_demux rsp_xbar_demux (
		.clk                (ddr2_afi_clk_clk),                    //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),       //          .channel
		.sink_data          (width_adapter_001_src_data),          //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),           //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),           //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),            //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),         //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),   //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)      //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (65),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (79),
		.IN_PKT_BYTE_CNT_L             (72),
		.IN_PKT_TRANS_COMPRESSED_READ  (66),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (80),
		.IN_PKT_BURST_SIZE_H           (83),
		.IN_PKT_BURST_SIZE_L           (81),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (71),
		.IN_PKT_BURST_TYPE_H           (85),
		.IN_PKT_BURST_TYPE_L           (84),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (317),
		.OUT_PKT_ADDR_L                (288),
		.OUT_PKT_DATA_H                (255),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (287),
		.OUT_PKT_BYTEEN_L              (256),
		.OUT_PKT_BYTE_CNT_H            (331),
		.OUT_PKT_BYTE_CNT_L            (324),
		.OUT_PKT_TRANS_COMPRESSED_READ (318),
		.OUT_PKT_BURST_SIZE_H          (335),
		.OUT_PKT_BURST_SIZE_L          (333),
		.OUT_PKT_RESPONSE_STATUS_H     (353),
		.OUT_PKT_RESPONSE_STATUS_L     (352),
		.OUT_PKT_TRANS_EXCLUSIVE       (323),
		.OUT_PKT_BURST_TYPE_H          (337),
		.OUT_PKT_BURST_TYPE_L          (336),
		.OUT_ST_DATA_W                 (354),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (ddr2_afi_clk_clk),                   //       clk.clk
		.reset                (rst_controller_002_reset_out_reset), // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src0_valid),          //      sink.valid
		.in_channel           (cmd_xbar_demux_src0_channel),        //          .channel
		.in_startofpacket     (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src0_endofpacket),    //          .endofpacket
		.in_ready             (cmd_xbar_demux_src0_ready),          //          .ready
		.in_data              (cmd_xbar_demux_src0_data),           //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (317),
		.IN_PKT_ADDR_L                 (288),
		.IN_PKT_DATA_H                 (255),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (287),
		.IN_PKT_BYTEEN_L               (256),
		.IN_PKT_BYTE_CNT_H             (331),
		.IN_PKT_BYTE_CNT_L             (324),
		.IN_PKT_TRANS_COMPRESSED_READ  (318),
		.IN_PKT_BURSTWRAP_H            (332),
		.IN_PKT_BURSTWRAP_L            (332),
		.IN_PKT_BURST_SIZE_H           (335),
		.IN_PKT_BURST_SIZE_L           (333),
		.IN_PKT_RESPONSE_STATUS_H      (353),
		.IN_PKT_RESPONSE_STATUS_L      (352),
		.IN_PKT_TRANS_EXCLUSIVE        (323),
		.IN_PKT_BURST_TYPE_H           (337),
		.IN_PKT_BURST_TYPE_L           (336),
		.IN_ST_DATA_W                  (354),
		.OUT_PKT_ADDR_H                (65),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (72),
		.OUT_PKT_TRANS_COMPRESSED_READ (66),
		.OUT_PKT_BURST_SIZE_H          (83),
		.OUT_PKT_BURST_SIZE_L          (81),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (71),
		.OUT_PKT_BURST_TYPE_H          (85),
		.OUT_PKT_BURST_TYPE_L          (84),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (ddr2_afi_clk_clk),                    //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_src_valid),                 //      sink.valid
		.in_channel           (id_router_src_channel),               //          .channel
		.in_startofpacket     (id_router_src_startofpacket),         //          .startofpacket
		.in_endofpacket       (id_router_src_endofpacket),           //          .endofpacket
		.in_ready             (id_router_src_ready),                 //          .ready
		.in_data              (id_router_src_data),                  //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

endmodule
